LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY sev_seg IS
PORT 	(bcd : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 neg : IN STD_LOGIC;
		 leds: OUT  STD_LOGIC_VECTOR(0 TO 6);
		 nleds: OUT  STD_LOGIC_VECTOR(0 TO 6));
	
END sev_seg;

ARCHITECTURE Behavior OF sev_seg IS
BEGIN
	PROCESS (bcd)
	BEGIN
		CASE bcd IS -- abcdefg
			WHEN "0000" => leds <= "1111110";--"0"
			WHEN "0001" => leds <= "0110000";--"1"
			WHEN "0010" => leds <= "1101101";--"2"
			WHEN "0011" => leds <= "1111001";--"3"
			WHEN "0100" => leds <= "0110011";--"4"
			WHEN "0101" => leds <= "1011011";--"5"
			WHEN "0110" => leds <= "1011111";--"6"
			WHEN "0111" => leds <= "1110000";--"7"
			WHEN "1000" => leds <= "1111111";--"8"
			WHEN "1001" => leds <= "1110011";--"9"
			WHEN "1010" => leds <= "1110111";--a
			WHEN "1011" => leds <= "0011111";--b
			WHEN "1100" => leds <= "1001110";--c
			WHEN "1101" => leds <= "0111101";--d
			WHEN "1110" => leds <= "1001111";--e
			WHEN "1111" => leds <= "1000111";--f
			WHEN OTHERS => leds <= "0000000";
END CASE;

END PROCESS;

PROCESS (Neg)
BEGIN
	CASE Neg IS
			WHEN '0' => nleds <= "0000000" ; --No negative sign
			WHEN '1' => nleds <= "0000001" ; --For negative sign
		END CASE;
	END PROCESS ;
END Behavior ;
                                           


